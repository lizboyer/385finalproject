[[0. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 5. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 5. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 5. 5. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 5. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 5. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 5. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 0. 5. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 0. 5. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 4. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 4. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 0. 1. 1. 0. 1. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 0. 0.
  0. 0. 0. 0. 0. 1. 0.]
 [0. 0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 0. 0. 4. 1.
  1. 1. 0. 0. 0. 0. 1.]
 [0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 0. 4. 4. 1. 1.
  1. 1. 0. 0. 0. 0. 0.]
 [0. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 5. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 0. 4. 1. 1. 1. 1.
  0. 1. 1. 0. 0. 0. 0.]
 [0. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 5. 5. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4.
  4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 1. 1. 1. 1.
  1. 1. 1. 1. 1. 1. 0.]
 [0. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 5. 5. 5. 5. 5. 0. 5. 5. 4. 4. 5. 4. 4.
  4. 4. 4. 4. 4. 5. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 1. 1. 1. 0. 1.
  1. 0. 1. 1. 1. 1. 0.]
 [0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 0. 0. 5. 5. 4. 5. 4. 4.
  4. 4. 4. 4. 4. 5. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 1. 1. 1. 1. 1.
  1. 1. 1. 0. 1. 1. 0.]
 [0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 0. 0. 0. 0. 5. 5. 5. 5. 4.
  4. 4. 4. 4. 4. 4. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 1. 0.
  1. 1. 1. 1. 1. 0. 0.]
 [0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 0. 0. 0. 0. 0. 5. 5. 4.
  4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 1. 1.
  1. 1. 1. 1. 1. 0. 0.]
 [4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 5. 0. 0. 0. 0. 5. 5. 5.
  4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 0. 0. 1. 1.
  1. 1. 1. 1. 0. 0. 0.]
 [4. 4. 4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 5. 5. 5. 0. 0. 5. 5. 5.
  5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 4. 4. 1. 1. 0. 0. 0. 1.
  1. 1. 1. 0. 0. 0. 0.]
 [4. 4. 0. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 0. 5. 5. 0. 5. 5. 5.
  5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 0. 4. 1. 1. 0. 0. 1. 1.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 5. 0. 5. 0. 5. 5. 5.
  5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 1. 1. 1. 1. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [4. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 5. 5. 5. 5. 0. 5. 0. 0. 0. 0.
  0. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]
 [0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 0. 4. 4. 0. 0. 0. 0. 0. 0. 0. 0. 0.
  0. 0. 0. 0. 0. 0. 0.]]
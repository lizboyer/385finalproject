
 module font_rom ( input [10:0]	addr, 
 output [7:0]	data 
); 
 
	parameter ADDR_WIDTH = 11; 
   parameter DATA_WIDTH =  8; 
	logic [ADDR_WIDTH-1:0] addr_reg; 
				 
	// ROM definition				 
	parameter [0:2**ADDR_WIDTH-1][DATA_WIDTH-1:0] ROM = [[7. 7. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 5. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 5. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 5. 5. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 5. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 5. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 5. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 7. 5. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 7. 5. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 7. 7. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 0. 0. 0. 0. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 0. 0. 0. 0. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 0. 0. 0. 0. 4. 4. 4. 0. 0. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 7. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 7. 7. 4. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 0. 4. 4. 4. 0. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 0. 0. 0. 0. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [7. 7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 0. 1. 1. 0. 1. 7. 7. 7. 7. 7. 7. 0. 0. 7.]
 [7. 7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 7. 7. 7. 7. 7. 0. 0. 1. 0.]
 [7. 7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 4. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 0. 0. 4. 1. 1. 1. 0. 0. 0. 0. 1.]
 [7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 0. 4. 4. 1. 1. 1. 1. 0. 0. 0. 0. 0.]
 [7. 4. 4. 4. 4. 4. 4. 4. 4. 4. 5. 5. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 0. 4. 1. 1. 1. 1. 0. 1. 1. 0. 0. 0. 7.]
 [7. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 5. 5. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 1. 1. 1. 1. 1. 1. 1. 1. 1. 1. 7.]
 [7. 4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 5. 5. 5. 5. 5. 7. 5. 5. 4. 4. 5. 4. 4. 4. 4. 4. 4. 4. 5. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 1. 1. 1. 0. 1. 1. 0. 1. 1. 1. 1. 7.]
 [7. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 7. 7. 5. 5. 4. 5. 4. 4. 4. 4. 4. 4. 4. 5. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 1. 1. 1. 1. 1. 1. 1. 1. 0. 1. 1. 7.]
 [7. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 7. 7. 7. 7. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 0. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 1. 0. 1. 1. 1. 1. 1. 7. 7.]
 [7. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 7. 7. 7. 7. 7. 5. 5. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 0. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 1. 1. 1. 1. 1. 1. 1. 1. 1. 7. 7.]
 [4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 5. 7. 7. 7. 7. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 0. 0. 0. 0. 0. 4. 4. 4. 1. 1. 0. 0. 1. 1. 1. 1. 1. 1. 7. 7. 7.]
 [4. 4. 4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 5. 5. 5. 7. 7. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 0. 7. 4. 4. 1. 1. 0. 0. 0. 1. 1. 1. 1. 7. 7. 7. 7.]
 [4. 4. 0. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 0. 5. 5. 7. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 4. 7. 7. 7. 4. 1. 1. 0. 0. 1. 1. 7. 7. 7. 7. 7. 7. 7.]
 [0. 0. 4. 4. 7. 7. 7. 7. 7. 7. 7. 7. 7. 5. 5. 5. 5. 5. 0. 5. 7. 5. 5. 5. 5. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 4. 7. 7. 7. 1. 1. 1. 1. 7. 7. 7. 7. 7. 7. 7. 7. 7.]
 [4. 4. 4. 7. 7. 7. 7. 7. 7. 7. 0. 0. 0. 0. 5. 5. 5. 5. 0. 5. 7. 7. 7. 0. 0. 5. 5. 4. 4. 4. 4. 4. 4. 4. 4. 4. 0. 4. 4. 7. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 7. 7. 7.]
 [0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 0. 4. 4. 4. 4. 4. 0. 4. 4. 7. 0. 0. 0. 0. 0. 0. 7. 7. 7. 7. 7. 7. 7. 7. 7.]]}; 
 
	assign data = ROM[addr]; 
 
 endmodule  